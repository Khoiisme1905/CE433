// system.v

// Generated using ACDS version 13.0sp1 232 at 2025.05.29.09:09:25

`timescale 1 ps / 1 ps
module system (
		input  wire       clk_clk,                          //                       clk.clk
		input  wire       reset_reset_n,                    //                     reset.reset_n
		input  wire [3:0] sw_in_external_connection_export, // sw_in_external_connection.export
		input  wire       sw_en_external_connection_export, // sw_en_external_connection.export
		output wire [6:0] hex_0_conduit_end_export,         //         hex_0_conduit_end.export
		output wire [6:0] hex_1_conduit_end_export          //         hex_1_conduit_end.export
	);

	wire         nios2_qsys_0_instruction_master_waitrequest;                                                         // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [16:0] nios2_qsys_0_instruction_master_address;                                                             // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire         nios2_qsys_0_instruction_master_read;                                                                // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                                            // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                                                                // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                                                  // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire  [16:0] nios2_qsys_0_data_master_address;                                                                    // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire         nios2_qsys_0_data_master_write;                                                                      // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire         nios2_qsys_0_data_master_read;                                                                       // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                                                   // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                                                                // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                                                 // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                           // nios2_qsys_0:jtag_debug_module_waitrequest -> nios2_qsys_0_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                             // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                               // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                 // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read;                                  // nios2_qsys_0_jtag_debug_module_translator:av_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                              // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                           // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                            // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                        // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire  [12:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                          // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                       // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                            // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                            // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                         // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire   [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                       // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire  [31:0] memory_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                    // Memory_0_avalon_slave_0_translator:av_writedata -> Memory_0:iData
	wire   [3:0] memory_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                      // Memory_0_avalon_slave_0_translator:av_address -> Memory_0:iAddress
	wire         memory_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                   // Memory_0_avalon_slave_0_translator:av_chipselect -> Memory_0:iChipSelect_n
	wire         memory_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                        // Memory_0_avalon_slave_0_translator:av_write -> Memory_0:iWrite_n
	wire         memory_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                         // Memory_0_avalon_slave_0_translator:av_read -> Memory_0:iRead_n
	wire  [31:0] memory_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                     // Memory_0:oData -> Memory_0_avalon_slave_0_translator:av_readdata
	wire   [7:0] hex_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                       // HEX_0_avalon_slave_0_translator:av_writedata -> HEX_0:iHex_Data
	wire         hex_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                      // HEX_0_avalon_slave_0_translator:av_chipselect -> HEX_0:iChip_select_n
	wire         hex_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                           // HEX_0_avalon_slave_0_translator:av_write -> HEX_0:iWrite_n
	wire  [31:0] fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                      // FMAX_0_avalon_slave_0_translator:av_writedata -> FMAX_0:iData
	wire   [1:0] fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                        // FMAX_0_avalon_slave_0_translator:av_address -> FMAX_0:iAddress
	wire         fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                     // FMAX_0_avalon_slave_0_translator:av_chipselect -> FMAX_0:iChipselect_n
	wire         fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                          // FMAX_0_avalon_slave_0_translator:av_write -> FMAX_0:iWrite_n
	wire         fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                           // FMAX_0_avalon_slave_0_translator:av_read -> FMAX_0:iRead_n
	wire  [31:0] fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                       // FMAX_0:oData -> FMAX_0_avalon_slave_0_translator:av_readdata
	wire   [7:0] hex_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                       // HEX_1_avalon_slave_0_translator:av_writedata -> HEX_1:iHex_Data
	wire         hex_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                      // HEX_1_avalon_slave_0_translator:av_chipselect -> HEX_1:iChip_select_n
	wire         hex_1_avalon_slave_0_translator_avalon_anti_slave_0_write;                                           // HEX_1_avalon_slave_0_translator:av_write -> HEX_1:iWrite_n
	wire   [1:0] sw_in_s1_translator_avalon_anti_slave_0_address;                                                     // SW_IN_s1_translator:av_address -> SW_IN:address
	wire  [31:0] sw_in_s1_translator_avalon_anti_slave_0_readdata;                                                    // SW_IN:readdata -> SW_IN_s1_translator:av_readdata
	wire   [1:0] sw_en_s1_translator_avalon_anti_slave_0_address;                                                     // SW_EN_s1_translator:av_address -> SW_EN:address
	wire  [31:0] sw_en_s1_translator_avalon_anti_slave_0_readdata;                                                    // SW_EN:readdata -> SW_EN_s1_translator:av_readdata
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                    // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                     // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                      // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [16:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                        // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                           // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                          // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                           // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                       // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                    // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                     // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                            // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                             // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [16:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                               // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                  // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                 // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                  // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                              // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                            // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire  [16:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [92:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [92:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire  [16:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [92:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [92:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [16:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [92:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [92:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // Memory_0_avalon_slave_0_translator:uav_waitrequest -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Memory_0_avalon_slave_0_translator:uav_burstcount
	wire  [31:0] memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                      // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Memory_0_avalon_slave_0_translator:uav_writedata
	wire  [16:0] memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                        // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Memory_0_avalon_slave_0_translator:uav_address
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                          // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Memory_0_avalon_slave_0_translator:uav_write
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                           // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Memory_0_avalon_slave_0_translator:uav_lock
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                           // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Memory_0_avalon_slave_0_translator:uav_read
	wire  [31:0] memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                       // Memory_0_avalon_slave_0_translator:uav_readdata -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // Memory_0_avalon_slave_0_translator:uav_readdatavalid -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Memory_0_avalon_slave_0_translator:uav_debugaccess
	wire   [3:0] memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Memory_0_avalon_slave_0_translator:uav_byteenable
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [92:0] memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                    // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [92:0] memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // HEX_0_avalon_slave_0_translator:uav_waitrequest -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [0:0] hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> HEX_0_avalon_slave_0_translator:uav_burstcount
	wire   [7:0] hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                         // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> HEX_0_avalon_slave_0_translator:uav_writedata
	wire  [16:0] hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                           // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> HEX_0_avalon_slave_0_translator:uav_address
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                             // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> HEX_0_avalon_slave_0_translator:uav_write
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                              // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> HEX_0_avalon_slave_0_translator:uav_lock
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                              // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> HEX_0_avalon_slave_0_translator:uav_read
	wire   [7:0] hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                          // HEX_0_avalon_slave_0_translator:uav_readdata -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // HEX_0_avalon_slave_0_translator:uav_readdatavalid -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> HEX_0_avalon_slave_0_translator:uav_debugaccess
	wire   [0:0] hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> HEX_0_avalon_slave_0_translator:uav_byteenable
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [65:0] hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                       // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [65:0] hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [9:0] hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // FMAX_0_avalon_slave_0_translator:uav_waitrequest -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> FMAX_0_avalon_slave_0_translator:uav_burstcount
	wire  [31:0] fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                        // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> FMAX_0_avalon_slave_0_translator:uav_writedata
	wire  [16:0] fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                          // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> FMAX_0_avalon_slave_0_translator:uav_address
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                            // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> FMAX_0_avalon_slave_0_translator:uav_write
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                             // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> FMAX_0_avalon_slave_0_translator:uav_lock
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                             // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> FMAX_0_avalon_slave_0_translator:uav_read
	wire  [31:0] fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                         // FMAX_0_avalon_slave_0_translator:uav_readdata -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // FMAX_0_avalon_slave_0_translator:uav_readdatavalid -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FMAX_0_avalon_slave_0_translator:uav_debugaccess
	wire   [3:0] fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> FMAX_0_avalon_slave_0_translator:uav_byteenable
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [92:0] fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                      // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [92:0] fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // HEX_1_avalon_slave_0_translator:uav_waitrequest -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [0:0] hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> HEX_1_avalon_slave_0_translator:uav_burstcount
	wire   [7:0] hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                         // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> HEX_1_avalon_slave_0_translator:uav_writedata
	wire  [16:0] hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                           // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> HEX_1_avalon_slave_0_translator:uav_address
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                             // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> HEX_1_avalon_slave_0_translator:uav_write
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                              // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> HEX_1_avalon_slave_0_translator:uav_lock
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                              // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> HEX_1_avalon_slave_0_translator:uav_read
	wire   [7:0] hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                          // HEX_1_avalon_slave_0_translator:uav_readdata -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // HEX_1_avalon_slave_0_translator:uav_readdatavalid -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> HEX_1_avalon_slave_0_translator:uav_debugaccess
	wire   [0:0] hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> HEX_1_avalon_slave_0_translator:uav_byteenable
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [65:0] hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                       // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [65:0] hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [9:0] hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // SW_IN_s1_translator:uav_waitrequest -> SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sw_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SW_IN_s1_translator:uav_burstcount
	wire  [31:0] sw_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SW_IN_s1_translator:uav_writedata
	wire  [16:0] sw_in_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_address -> SW_IN_s1_translator:uav_address
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_write -> SW_IN_s1_translator:uav_write
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SW_IN_s1_translator:uav_lock
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_read -> SW_IN_s1_translator:uav_read
	wire  [31:0] sw_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // SW_IN_s1_translator:uav_readdata -> SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // SW_IN_s1_translator:uav_readdatavalid -> SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SW_IN_s1_translator:uav_debugaccess
	wire   [3:0] sw_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // SW_IN_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SW_IN_s1_translator:uav_byteenable
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [92:0] sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [92:0] sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // SW_IN_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // SW_IN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SW_IN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sw_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // SW_IN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SW_IN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // SW_IN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SW_IN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // SW_EN_s1_translator:uav_waitrequest -> SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sw_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SW_EN_s1_translator:uav_burstcount
	wire  [31:0] sw_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SW_EN_s1_translator:uav_writedata
	wire  [16:0] sw_en_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_address -> SW_EN_s1_translator:uav_address
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_write -> SW_EN_s1_translator:uav_write
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SW_EN_s1_translator:uav_lock
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_read -> SW_EN_s1_translator:uav_read
	wire  [31:0] sw_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // SW_EN_s1_translator:uav_readdata -> SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // SW_EN_s1_translator:uav_readdatavalid -> SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SW_EN_s1_translator:uav_debugaccess
	wire   [3:0] sw_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // SW_EN_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SW_EN_s1_translator:uav_byteenable
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [92:0] sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [92:0] sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // SW_EN_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // SW_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SW_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sw_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // SW_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SW_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // SW_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SW_EN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                 // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [91:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [91:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [91:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [91:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_001:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [91:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_002:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                          // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [91:0] memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                           // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_003:sink_ready -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                             // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [64:0] hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                              // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_004:sink_ready -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                            // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [91:0] fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                             // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_005:sink_ready -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                             // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [64:0] hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                              // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_006:sink_ready -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // SW_IN_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // SW_IN_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // SW_IN_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [91:0] sw_in_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // SW_IN_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         sw_in_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_007:sink_ready -> SW_IN_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // SW_EN_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // SW_EN_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // SW_EN_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [91:0] sw_en_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // SW_EN_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         sw_en_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_008:sink_ready -> SW_EN_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         burst_adapter_source0_endofpacket;                                                                   // burst_adapter:source0_endofpacket -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                         // burst_adapter:source0_valid -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                                 // burst_adapter:source0_startofpacket -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [64:0] burst_adapter_source0_data;                                                                          // burst_adapter:source0_data -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                         // HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [8:0] burst_adapter_source0_channel;                                                                       // burst_adapter:source0_channel -> HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_001_source0_endofpacket;                                                               // burst_adapter_001:source0_endofpacket -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_001_source0_valid;                                                                     // burst_adapter_001:source0_valid -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_001_source0_startofpacket;                                                             // burst_adapter_001:source0_startofpacket -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [64:0] burst_adapter_001_source0_data;                                                                      // burst_adapter_001:source0_data -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_001_source0_ready;                                                                     // HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [8:0] burst_adapter_001_source0_channel;                                                                   // burst_adapter_001:source0_channel -> HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                      // rst_controller:reset_out -> [FMAX_0:iReset_n, FMAX_0_avalon_slave_0_translator:reset, FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, HEX_0:iReset_n, HEX_0_avalon_slave_0_translator:reset, HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, HEX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, HEX_1:iReset_n, HEX_1_avalon_slave_0_translator:reset, HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, HEX_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Memory_0:iReset_n, Memory_0_avalon_slave_0_translator:reset, Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire         rst_controller_reset_out_reset_req;                                                                  // rst_controller:reset_req -> onchip_memory2_0:reset_req
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                                                          // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                                                  // rst_controller_001:reset_out -> [SW_EN:reset_n, SW_EN_s1_translator:reset, SW_EN_s1_translator_avalon_universal_slave_0_agent:reset, SW_EN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SW_IN:reset_n, SW_IN_s1_translator:reset, SW_IN_s1_translator_avalon_universal_slave_0_agent:reset, SW_IN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_007:reset, id_router_008:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                     // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                           // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                   // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [91:0] cmd_xbar_demux_src0_data;                                                                            // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [8:0] cmd_xbar_demux_src0_channel;                                                                         // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                           // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                     // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                           // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                   // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [91:0] cmd_xbar_demux_src1_data;                                                                            // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [8:0] cmd_xbar_demux_src1_channel;                                                                         // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                           // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                     // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                           // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                   // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [91:0] cmd_xbar_demux_src2_data;                                                                            // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [8:0] cmd_xbar_demux_src2_channel;                                                                         // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                           // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                     // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                           // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                   // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [91:0] cmd_xbar_demux_src3_data;                                                                            // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [8:0] cmd_xbar_demux_src3_channel;                                                                         // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                           // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_src4_endofpacket;                                                                     // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                           // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                   // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [91:0] cmd_xbar_demux_src4_data;                                                                            // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire   [8:0] cmd_xbar_demux_src4_channel;                                                                         // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire         cmd_xbar_demux_src4_ready;                                                                           // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire         cmd_xbar_demux_src5_endofpacket;                                                                     // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                                           // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                                   // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [91:0] cmd_xbar_demux_src5_data;                                                                            // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [8:0] cmd_xbar_demux_src5_channel;                                                                         // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire         cmd_xbar_demux_src5_ready;                                                                           // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire         cmd_xbar_demux_src6_endofpacket;                                                                     // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                                           // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                                   // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [91:0] cmd_xbar_demux_src6_data;                                                                            // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire   [8:0] cmd_xbar_demux_src6_channel;                                                                         // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire         cmd_xbar_demux_src6_ready;                                                                           // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                 // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                       // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                               // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [91:0] cmd_xbar_demux_001_src0_data;                                                                        // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src0_channel;                                                                     // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                       // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                 // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                       // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                               // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [91:0] cmd_xbar_demux_001_src1_data;                                                                        // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src1_channel;                                                                     // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                       // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                 // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                       // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                               // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [91:0] cmd_xbar_demux_001_src2_data;                                                                        // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src2_channel;                                                                     // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                       // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                 // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                       // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                               // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [91:0] cmd_xbar_demux_001_src3_data;                                                                        // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src3_channel;                                                                     // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                       // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                 // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                       // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                               // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [91:0] cmd_xbar_demux_001_src4_data;                                                                        // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src4_channel;                                                                     // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire         cmd_xbar_demux_001_src4_ready;                                                                       // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                 // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                       // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                               // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [91:0] cmd_xbar_demux_001_src5_data;                                                                        // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src5_channel;                                                                     // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	wire         cmd_xbar_demux_001_src5_ready;                                                                       // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                 // cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                       // cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                               // cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [91:0] cmd_xbar_demux_001_src6_data;                                                                        // cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	wire   [8:0] cmd_xbar_demux_001_src6_channel;                                                                     // cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	wire         cmd_xbar_demux_001_src6_ready;                                                                       // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                 // cmd_xbar_demux_001:src7_endofpacket -> SW_IN_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                       // cmd_xbar_demux_001:src7_valid -> SW_IN_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                               // cmd_xbar_demux_001:src7_startofpacket -> SW_IN_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [91:0] cmd_xbar_demux_001_src7_data;                                                                        // cmd_xbar_demux_001:src7_data -> SW_IN_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src7_channel;                                                                     // cmd_xbar_demux_001:src7_channel -> SW_IN_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                 // cmd_xbar_demux_001:src8_endofpacket -> SW_EN_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                       // cmd_xbar_demux_001:src8_valid -> SW_EN_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                               // cmd_xbar_demux_001:src8_startofpacket -> SW_EN_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [91:0] cmd_xbar_demux_001_src8_data;                                                                        // cmd_xbar_demux_001:src8_data -> SW_EN_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_demux_001_src8_channel;                                                                     // cmd_xbar_demux_001:src8_channel -> SW_EN_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                     // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                           // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                   // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [91:0] rsp_xbar_demux_src0_data;                                                                            // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [8:0] rsp_xbar_demux_src0_channel;                                                                         // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                           // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                     // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                           // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                   // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [91:0] rsp_xbar_demux_src1_data;                                                                            // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [8:0] rsp_xbar_demux_src1_channel;                                                                         // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                           // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                 // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                       // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                               // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [91:0] rsp_xbar_demux_001_src0_data;                                                                        // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src0_channel;                                                                     // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                       // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                 // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                       // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                               // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [91:0] rsp_xbar_demux_001_src1_data;                                                                        // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [8:0] rsp_xbar_demux_001_src1_channel;                                                                     // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                       // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                 // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                       // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                               // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [91:0] rsp_xbar_demux_002_src0_data;                                                                        // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [8:0] rsp_xbar_demux_002_src0_channel;                                                                     // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                       // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                 // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                       // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                               // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [91:0] rsp_xbar_demux_002_src1_data;                                                                        // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [8:0] rsp_xbar_demux_002_src1_channel;                                                                     // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                       // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                 // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                       // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                               // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [91:0] rsp_xbar_demux_003_src0_data;                                                                        // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [8:0] rsp_xbar_demux_003_src0_channel;                                                                     // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                       // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                                 // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                       // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                               // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [91:0] rsp_xbar_demux_003_src1_data;                                                                        // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [8:0] rsp_xbar_demux_003_src1_channel;                                                                     // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                       // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                 // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                       // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                               // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [91:0] rsp_xbar_demux_004_src0_data;                                                                        // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [8:0] rsp_xbar_demux_004_src0_channel;                                                                     // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                       // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_004_src1_endofpacket;                                                                 // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src1_valid;                                                                       // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src1_startofpacket;                                                               // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [91:0] rsp_xbar_demux_004_src1_data;                                                                        // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [8:0] rsp_xbar_demux_004_src1_channel;                                                                     // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src1_ready;                                                                       // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                 // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                       // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                               // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [91:0] rsp_xbar_demux_005_src0_data;                                                                        // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [8:0] rsp_xbar_demux_005_src0_channel;                                                                     // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                       // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_005_src1_endofpacket;                                                                 // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src1_valid;                                                                       // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src1_startofpacket;                                                               // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [91:0] rsp_xbar_demux_005_src1_data;                                                                        // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	wire   [8:0] rsp_xbar_demux_005_src1_channel;                                                                     // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src1_ready;                                                                       // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                 // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                       // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                               // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [91:0] rsp_xbar_demux_006_src0_data;                                                                        // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire   [8:0] rsp_xbar_demux_006_src0_channel;                                                                     // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                       // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_006_src1_endofpacket;                                                                 // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src1_valid;                                                                       // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src1_startofpacket;                                                               // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [91:0] rsp_xbar_demux_006_src1_data;                                                                        // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	wire   [8:0] rsp_xbar_demux_006_src1_channel;                                                                     // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src1_ready;                                                                       // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                 // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                       // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                               // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [91:0] rsp_xbar_demux_007_src0_data;                                                                        // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [8:0] rsp_xbar_demux_007_src0_channel;                                                                     // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                       // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                 // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                       // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                               // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [91:0] rsp_xbar_demux_008_src0_data;                                                                        // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [8:0] rsp_xbar_demux_008_src0_channel;                                                                     // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                       // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         addr_router_src_endofpacket;                                                                         // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                               // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                       // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [91:0] addr_router_src_data;                                                                                // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [8:0] addr_router_src_channel;                                                                             // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                               // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                        // rsp_xbar_mux:src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                              // rsp_xbar_mux:src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                      // rsp_xbar_mux:src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [91:0] rsp_xbar_mux_src_data;                                                                               // rsp_xbar_mux:src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] rsp_xbar_mux_src_channel;                                                                            // rsp_xbar_mux:src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                              // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                     // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                           // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                   // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [91:0] addr_router_001_src_data;                                                                            // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [8:0] addr_router_001_src_channel;                                                                         // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                           // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                    // rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                          // rsp_xbar_mux_001:src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                  // rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [91:0] rsp_xbar_mux_001_src_data;                                                                           // rsp_xbar_mux_001:src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [8:0] rsp_xbar_mux_001_src_channel;                                                                        // rsp_xbar_mux_001:src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                          // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                        // cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                              // cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                      // cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [91:0] cmd_xbar_mux_src_data;                                                                               // cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_src_channel;                                                                            // cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                           // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                 // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                         // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [91:0] id_router_src_data;                                                                                  // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [8:0] id_router_src_channel;                                                                               // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                 // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                    // cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                          // cmd_xbar_mux_001:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                  // cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [91:0] cmd_xbar_mux_001_src_data;                                                                           // cmd_xbar_mux_001:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_001_src_channel;                                                                        // cmd_xbar_mux_001:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                       // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                             // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                     // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [91:0] id_router_001_src_data;                                                                              // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [8:0] id_router_001_src_channel;                                                                           // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                             // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                    // cmd_xbar_mux_002:src_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                          // cmd_xbar_mux_002:src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                  // cmd_xbar_mux_002:src_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [91:0] cmd_xbar_mux_002_src_data;                                                                           // cmd_xbar_mux_002:src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_002_src_channel;                                                                        // cmd_xbar_mux_002:src_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                       // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                             // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                     // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [91:0] id_router_002_src_data;                                                                              // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [8:0] id_router_002_src_channel;                                                                           // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                             // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                    // cmd_xbar_mux_003:src_endofpacket -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                          // cmd_xbar_mux_003:src_valid -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                                  // cmd_xbar_mux_003:src_startofpacket -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [91:0] cmd_xbar_mux_003_src_data;                                                                           // cmd_xbar_mux_003:src_data -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_003_src_channel;                                                                        // cmd_xbar_mux_003:src_channel -> Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                          // Memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire         id_router_003_src_endofpacket;                                                                       // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                             // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                     // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [91:0] id_router_003_src_data;                                                                              // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [8:0] id_router_003_src_channel;                                                                           // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                             // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_mux_005_src_endofpacket;                                                                    // cmd_xbar_mux_005:src_endofpacket -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_005_src_valid;                                                                          // cmd_xbar_mux_005:src_valid -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_005_src_startofpacket;                                                                  // cmd_xbar_mux_005:src_startofpacket -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [91:0] cmd_xbar_mux_005_src_data;                                                                           // cmd_xbar_mux_005:src_data -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [8:0] cmd_xbar_mux_005_src_channel;                                                                        // cmd_xbar_mux_005:src_channel -> FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_005_src_ready;                                                                          // FMAX_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire         id_router_005_src_endofpacket;                                                                       // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                             // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                     // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [91:0] id_router_005_src_data;                                                                              // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [8:0] id_router_005_src_channel;                                                                           // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                             // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                       // SW_IN_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                       // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                             // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                     // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [91:0] id_router_007_src_data;                                                                              // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [8:0] id_router_007_src_channel;                                                                           // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                             // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                       // SW_EN_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                       // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                             // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                     // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [91:0] id_router_008_src_data;                                                                              // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [8:0] id_router_008_src_channel;                                                                           // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                             // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_mux_004_src_endofpacket;                                                                    // cmd_xbar_mux_004:src_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_mux_004_src_valid;                                                                          // cmd_xbar_mux_004:src_valid -> width_adapter:in_valid
	wire         cmd_xbar_mux_004_src_startofpacket;                                                                  // cmd_xbar_mux_004:src_startofpacket -> width_adapter:in_startofpacket
	wire  [91:0] cmd_xbar_mux_004_src_data;                                                                           // cmd_xbar_mux_004:src_data -> width_adapter:in_data
	wire   [8:0] cmd_xbar_mux_004_src_channel;                                                                        // cmd_xbar_mux_004:src_channel -> width_adapter:in_channel
	wire         cmd_xbar_mux_004_src_ready;                                                                          // width_adapter:in_ready -> cmd_xbar_mux_004:src_ready
	wire         width_adapter_src_endofpacket;                                                                       // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                             // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                     // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [64:0] width_adapter_src_data;                                                                              // width_adapter:out_data -> burst_adapter:sink0_data
	wire         width_adapter_src_ready;                                                                             // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [8:0] width_adapter_src_channel;                                                                           // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire         id_router_004_src_endofpacket;                                                                       // id_router_004:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_004_src_valid;                                                                             // id_router_004:src_valid -> width_adapter_001:in_valid
	wire         id_router_004_src_startofpacket;                                                                     // id_router_004:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [64:0] id_router_004_src_data;                                                                              // id_router_004:src_data -> width_adapter_001:in_data
	wire   [8:0] id_router_004_src_channel;                                                                           // id_router_004:src_channel -> width_adapter_001:in_channel
	wire         id_router_004_src_ready;                                                                             // width_adapter_001:in_ready -> id_router_004:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                   // width_adapter_001:out_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                         // width_adapter_001:out_valid -> rsp_xbar_demux_004:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                                 // width_adapter_001:out_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [91:0] width_adapter_001_src_data;                                                                          // width_adapter_001:out_data -> rsp_xbar_demux_004:sink_data
	wire         width_adapter_001_src_ready;                                                                         // rsp_xbar_demux_004:sink_ready -> width_adapter_001:out_ready
	wire   [8:0] width_adapter_001_src_channel;                                                                       // width_adapter_001:out_channel -> rsp_xbar_demux_004:sink_channel
	wire         cmd_xbar_mux_006_src_endofpacket;                                                                    // cmd_xbar_mux_006:src_endofpacket -> width_adapter_002:in_endofpacket
	wire         cmd_xbar_mux_006_src_valid;                                                                          // cmd_xbar_mux_006:src_valid -> width_adapter_002:in_valid
	wire         cmd_xbar_mux_006_src_startofpacket;                                                                  // cmd_xbar_mux_006:src_startofpacket -> width_adapter_002:in_startofpacket
	wire  [91:0] cmd_xbar_mux_006_src_data;                                                                           // cmd_xbar_mux_006:src_data -> width_adapter_002:in_data
	wire   [8:0] cmd_xbar_mux_006_src_channel;                                                                        // cmd_xbar_mux_006:src_channel -> width_adapter_002:in_channel
	wire         cmd_xbar_mux_006_src_ready;                                                                          // width_adapter_002:in_ready -> cmd_xbar_mux_006:src_ready
	wire         width_adapter_002_src_endofpacket;                                                                   // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire         width_adapter_002_src_valid;                                                                         // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire         width_adapter_002_src_startofpacket;                                                                 // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [64:0] width_adapter_002_src_data;                                                                          // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire         width_adapter_002_src_ready;                                                                         // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire   [8:0] width_adapter_002_src_channel;                                                                       // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire         id_router_006_src_endofpacket;                                                                       // id_router_006:src_endofpacket -> width_adapter_003:in_endofpacket
	wire         id_router_006_src_valid;                                                                             // id_router_006:src_valid -> width_adapter_003:in_valid
	wire         id_router_006_src_startofpacket;                                                                     // id_router_006:src_startofpacket -> width_adapter_003:in_startofpacket
	wire  [64:0] id_router_006_src_data;                                                                              // id_router_006:src_data -> width_adapter_003:in_data
	wire   [8:0] id_router_006_src_channel;                                                                           // id_router_006:src_channel -> width_adapter_003:in_channel
	wire         id_router_006_src_ready;                                                                             // width_adapter_003:in_ready -> id_router_006:src_ready
	wire         width_adapter_003_src_endofpacket;                                                                   // width_adapter_003:out_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         width_adapter_003_src_valid;                                                                         // width_adapter_003:out_valid -> rsp_xbar_demux_006:sink_valid
	wire         width_adapter_003_src_startofpacket;                                                                 // width_adapter_003:out_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [91:0] width_adapter_003_src_data;                                                                          // width_adapter_003:out_data -> rsp_xbar_demux_006:sink_data
	wire         width_adapter_003_src_ready;                                                                         // rsp_xbar_demux_006:sink_ready -> width_adapter_003:out_ready
	wire   [8:0] width_adapter_003_src_channel;                                                                       // width_adapter_003:out_channel -> rsp_xbar_demux_006:sink_channel
	wire         irq_mapper_receiver0_irq;                                                                            // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                                                              // irq_mapper:sender_irq -> nios2_qsys_0:d_irq

	system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                                   //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                           //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                                       //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                             //       .reset_req
	);

	system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	Memory #(
		.DATA_WIDTH    (32),
		.ADDRESS_WIDTH (4)
	) memory_0 (
		.iRead_n       (~memory_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read_n
		.iWrite_n      (~memory_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write_n
		.iAddress      (memory_0_avalon_slave_0_translator_avalon_anti_slave_0_address),     //               .address
		.iData         (memory_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //               .writedata
		.oData         (memory_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //               .readdata
		.iChipSelect_n (~memory_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect_n
		.iClk          (clk_clk),                                                            //     clock_sink.clk
		.iReset_n      (~rst_controller_reset_out_reset)                                     //     reset_sink.reset_n
	);

	MAX_IP fmax_0 (
		.iChipselect_n (~fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), // avalon_slave_0.chipselect_n
		.iWrite_n      (~fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write_n
		.iRead_n       (~fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //               .read_n
		.iAddress      (fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_address),     //               .address
		.iData         (fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //               .writedata
		.oData         (fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //               .readdata
		.iClk          (clk_clk),                                                          //     clock_sink.clk
		.iReset_n      (~rst_controller_reset_out_reset)                                   //     reset_sink.reset_n
	);

	HEX_Control hex_0 (
		.iWrite_n       (~hex_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      // avalon_slave_0.write_n
		.iHex_Data      (hex_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //               .writedata
		.iChip_select_n (~hex_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect_n
		.iClk           (clk_clk),                                                         //     clock_sink.clk
		.iReset_n       (~rst_controller_reset_out_reset),                                 //     reset_sink.reset_n
		.oHex_Display   (hex_0_conduit_end_export)                                         //    conduit_end.export
	);

	system_SW_IN sw_in (
		.clk      (clk_clk),                                          //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address  (sw_in_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (sw_in_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (sw_in_external_connection_export)                  // external_connection.export
	);

	system_SW_EN sw_en (
		.clk      (clk_clk),                                          //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address  (sw_en_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (sw_en_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (sw_en_external_connection_export)                  // external_connection.export
	);

	HEX_Control hex_1 (
		.iWrite_n       (~hex_1_avalon_slave_0_translator_avalon_anti_slave_0_write),      // avalon_slave_0.write_n
		.iHex_Data      (hex_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //               .writedata
		.iChip_select_n (~hex_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect_n
		.iClk           (clk_clk),                                                         //     clock_sink.clk
		.iReset_n       (~rst_controller_reset_out_reset),                                 //     reset_sink.reset_n
		.oHex_Display   (hex_1_conduit_end_export)                                         //    conduit_end.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (17),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (17),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                      (clk_clk),                                                                            //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                               //               (terminated)
		.av_byteenable            (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                                               //               (terminated)
		.av_readdatavalid         (),                                                                                   //               (terminated)
		.av_write                 (1'b0),                                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock                  (1'b0),                                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                                               //               (terminated)
		.uav_clken                (),                                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                                               //               (terminated)
		.uav_response             (2'b00),                                                                              //               (terminated)
		.av_response              (),                                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (17),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (17),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2_qsys_0_data_master_translator (
		.clk                      (clk_clk),                                                                     //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata             (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) memory_0_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (memory_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (memory_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (memory_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (memory_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (memory_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (memory_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_byteenable            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_debugaccess           (),                                                                                   //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex_0_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address              (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (hex_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (hex_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                                //              (terminated)
		.av_read                  (),                                                                                //              (terminated)
		.av_readdata              (8'b10101101),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                //              (terminated)
		.av_burstcount            (),                                                                                //              (terminated)
		.av_byteenable            (),                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                //              (terminated)
		.av_lock                  (),                                                                                //              (terminated)
		.av_clken                 (),                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                //              (terminated)
		.uav_response             (),                                                                                //              (terminated)
		.av_response              (2'b00),                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fmax_0_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (fmax_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_byteenable            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex_1_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address              (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (hex_1_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (hex_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                                //              (terminated)
		.av_read                  (),                                                                                //              (terminated)
		.av_readdata              (8'b10101101),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                //              (terminated)
		.av_burstcount            (),                                                                                //              (terminated)
		.av_byteenable            (),                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                //              (terminated)
		.av_lock                  (),                                                                                //              (terminated)
		.av_clken                 (),                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                //              (terminated)
		.uav_response             (),                                                                                //              (terminated)
		.av_response              (2'b00),                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sw_in_s1_translator (
		.clk                      (clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sw_in_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sw_in_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                    //              (terminated)
		.av_read                  (),                                                                    //              (terminated)
		.av_writedata             (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_chipselect            (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sw_en_s1_translator (
		.clk                      (clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sw_en_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sw_en_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                    //              (terminated)
		.av_read                  (),                                                                    //              (terminated)
		.av_writedata             (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_chipselect            (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.PKT_BURST_TYPE_H          (69),
		.PKT_BURST_TYPE_L          (68),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_TRANS_EXCLUSIVE       (58),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (82),
		.PKT_THREAD_ID_L           (82),
		.PKT_CACHE_H               (89),
		.PKT_CACHE_L               (86),
		.PKT_DATA_SIDEBAND_H       (71),
		.PKT_DATA_SIDEBAND_L       (71),
		.PKT_QOS_H                 (73),
		.PKT_QOS_L                 (73),
		.PKT_ADDR_SIDEBAND_H       (70),
		.PKT_ADDR_SIDEBAND_L       (70),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.ST_DATA_W                 (92),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                     //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                      //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                       //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                                //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                      //          .ready
		.av_response             (),                                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.PKT_BURST_TYPE_H          (69),
		.PKT_BURST_TYPE_L          (68),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_TRANS_EXCLUSIVE       (58),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (78),
		.PKT_THREAD_ID_H           (82),
		.PKT_THREAD_ID_L           (82),
		.PKT_CACHE_H               (89),
		.PKT_CACHE_L               (86),
		.PKT_DATA_SIDEBAND_H       (71),
		.PKT_DATA_SIDEBAND_L       (71),
		.PKT_QOS_H                 (73),
		.PKT_QOS_L                 (73),
		.PKT_ADDR_SIDEBAND_H       (70),
		.PKT_ADDR_SIDEBAND_L       (70),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.ST_DATA_W                 (92),
		.ST_CHANNEL_W              (9),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                              //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                           //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                            //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                         //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                                     //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                           //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (92),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (93),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (92),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (93),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (92),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                       //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (93),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (92),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                                 //                .channel
		.rf_sink_ready           (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (93),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (45),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (25),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (26),
		.PKT_TRANS_POSTED          (27),
		.PKT_TRANS_WRITE           (28),
		.PKT_TRANS_READ            (29),
		.PKT_TRANS_LOCK            (30),
		.PKT_SRC_ID_H              (50),
		.PKT_SRC_ID_L              (47),
		.PKT_DEST_ID_H             (54),
		.PKT_DEST_ID_L             (51),
		.PKT_BURSTWRAP_H           (37),
		.PKT_BURSTWRAP_L           (35),
		.PKT_BYTE_CNT_H            (34),
		.PKT_BYTE_CNT_L            (32),
		.PKT_PROTECTION_H          (58),
		.PKT_PROTECTION_L          (56),
		.PKT_RESPONSE_STATUS_H     (64),
		.PKT_RESPONSE_STATUS_L     (63),
		.PKT_BURST_SIZE_H          (40),
		.PKT_BURST_SIZE_L          (38),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (65),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                               //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                               //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                         //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                             //                .channel
		.rf_sink_ready           (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (66),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (92),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                               //                .channel
		.rf_sink_ready           (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (93),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (45),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (25),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (26),
		.PKT_TRANS_POSTED          (27),
		.PKT_TRANS_WRITE           (28),
		.PKT_TRANS_READ            (29),
		.PKT_TRANS_LOCK            (30),
		.PKT_SRC_ID_H              (50),
		.PKT_SRC_ID_L              (47),
		.PKT_DEST_ID_H             (54),
		.PKT_DEST_ID_L             (51),
		.PKT_BURSTWRAP_H           (37),
		.PKT_BURSTWRAP_L           (35),
		.PKT_BYTE_CNT_H            (34),
		.PKT_BYTE_CNT_L            (32),
		.PKT_PROTECTION_H          (58),
		.PKT_PROTECTION_L          (56),
		.PKT_RESPONSE_STATUS_H     (64),
		.PKT_RESPONSE_STATUS_L     (63),
		.PKT_BURST_SIZE_H          (40),
		.PKT_BURST_SIZE_L          (38),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (65),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                           //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                           //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                            //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                     //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                         //                .channel
		.rf_sink_ready           (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (66),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (92),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sw_in_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sw_in_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                               //                .channel
		.rf_sink_ready           (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sw_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sw_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sw_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sw_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sw_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sw_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (93),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sw_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sw_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (9),
		.ST_DATA_W                 (92),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sw_en_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sw_en_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                               //                .channel
		.rf_sink_ready           (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sw_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sw_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sw_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sw_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sw_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sw_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (93),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sw_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sw_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	system_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	system_id_router id_router (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	system_id_router id_router_001 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                        //       src.ready
		.src_valid          (id_router_001_src_valid),                                                        //          .valid
		.src_data           (id_router_001_src_data),                                                         //          .data
		.src_channel        (id_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	system_id_router id_router_002 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                  //          .valid
		.src_data           (id_router_002_src_data),                                                                   //          .data
		.src_channel        (id_router_002_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                             //          .endofpacket
	);

	system_id_router id_router_003 (
		.sink_ready         (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (memory_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                            //       src.ready
		.src_valid          (id_router_003_src_valid),                                                            //          .valid
		.src_data           (id_router_003_src_data),                                                             //          .data
		.src_channel        (id_router_003_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                       //          .endofpacket
	);

	system_id_router_004 id_router_004 (
		.sink_ready         (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                         //       src.ready
		.src_valid          (id_router_004_src_valid),                                                         //          .valid
		.src_data           (id_router_004_src_data),                                                          //          .data
		.src_channel        (id_router_004_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                    //          .endofpacket
	);

	system_id_router id_router_005 (
		.sink_ready         (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fmax_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                          //       src.ready
		.src_valid          (id_router_005_src_valid),                                                          //          .valid
		.src_data           (id_router_005_src_data),                                                           //          .data
		.src_channel        (id_router_005_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                     //          .endofpacket
	);

	system_id_router_004 id_router_006 (
		.sink_ready         (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                         //       src.ready
		.src_valid          (id_router_006_src_valid),                                                         //          .valid
		.src_data           (id_router_006_src_data),                                                          //          .data
		.src_channel        (id_router_006_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                    //          .endofpacket
	);

	system_id_router_007 id_router_007 (
		.sink_ready         (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sw_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                             //       src.ready
		.src_valid          (id_router_007_src_valid),                                             //          .valid
		.src_data           (id_router_007_src_data),                                              //          .data
		.src_channel        (id_router_007_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                        //          .endofpacket
	);

	system_id_router_007 id_router_008 (
		.sink_ready         (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sw_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                             //       src.ready
		.src_valid          (id_router_008_src_valid),                                             //          .valid
		.src_data           (id_router_008_src_data),                                              //          .data
		.src_channel        (id_router_008_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                        //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (25),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (45),
		.PKT_BYTE_CNT_H            (34),
		.PKT_BYTE_CNT_L            (32),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (40),
		.PKT_BURST_SIZE_L          (38),
		.PKT_BURST_TYPE_H          (42),
		.PKT_BURST_TYPE_L          (41),
		.PKT_BURSTWRAP_H           (37),
		.PKT_BURSTWRAP_L           (35),
		.PKT_TRANS_COMPRESSED_READ (26),
		.PKT_TRANS_WRITE           (28),
		.PKT_TRANS_READ            (29),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (65),
		.ST_CHANNEL_W              (9),
		.OUT_BYTE_CNT_H            (32),
		.OUT_BURSTWRAP_H           (37),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clk_clk),                             //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (25),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (45),
		.PKT_BYTE_CNT_H            (34),
		.PKT_BYTE_CNT_L            (32),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (40),
		.PKT_BURST_SIZE_L          (38),
		.PKT_BURST_TYPE_H          (42),
		.PKT_BURST_TYPE_L          (41),
		.PKT_BURSTWRAP_H           (37),
		.PKT_BURSTWRAP_L           (35),
		.PKT_TRANS_COMPRESSED_READ (26),
		.PKT_TRANS_WRITE           (28),
		.PKT_TRANS_READ            (29),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (65),
		.ST_CHANNEL_W              (9),
		.OUT_BYTE_CNT_H            (32),
		.OUT_BURSTWRAP_H           (37),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                    //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket),   //          .endofpacket
		.src6_ready         (cmd_xbar_demux_src6_ready),         //      src6.ready
		.src6_valid         (cmd_xbar_demux_src6_valid),         //          .valid
		.src6_data          (cmd_xbar_demux_src6_data),          //          .data
		.src6_channel       (cmd_xbar_demux_src6_channel),       //          .channel
		.src6_startofpacket (cmd_xbar_demux_src6_startofpacket), //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_src6_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //      src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //      src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.src8_ready         (cmd_xbar_demux_001_src8_ready),         //      src8.ready
		.src8_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.src8_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.src8_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.src8_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_mux cmd_xbar_mux_006 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src6_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src6_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux_007 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux_007 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src1_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src1_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (52),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (61),
		.IN_PKT_BYTE_CNT_L             (59),
		.IN_PKT_TRANS_COMPRESSED_READ  (53),
		.IN_PKT_BURSTWRAP_H            (64),
		.IN_PKT_BURSTWRAP_L            (62),
		.IN_PKT_BURST_SIZE_H           (67),
		.IN_PKT_BURST_SIZE_L           (65),
		.IN_PKT_RESPONSE_STATUS_H      (91),
		.IN_PKT_RESPONSE_STATUS_L      (90),
		.IN_PKT_TRANS_EXCLUSIVE        (58),
		.IN_PKT_BURST_TYPE_H           (69),
		.IN_PKT_BURST_TYPE_L           (68),
		.IN_ST_DATA_W                  (92),
		.OUT_PKT_ADDR_H                (25),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (34),
		.OUT_PKT_BYTE_CNT_L            (32),
		.OUT_PKT_TRANS_COMPRESSED_READ (26),
		.OUT_PKT_BURST_SIZE_H          (40),
		.OUT_PKT_BURST_SIZE_L          (38),
		.OUT_PKT_RESPONSE_STATUS_H     (64),
		.OUT_PKT_RESPONSE_STATUS_L     (63),
		.OUT_PKT_TRANS_EXCLUSIVE       (31),
		.OUT_PKT_BURST_TYPE_H          (42),
		.OUT_PKT_BURST_TYPE_L          (41),
		.OUT_ST_DATA_W                 (65),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clk_clk),                            //       clk.clk
		.reset                (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_mux_004_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_004_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_004_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_004_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_004_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_004_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (25),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (34),
		.IN_PKT_BYTE_CNT_L             (32),
		.IN_PKT_TRANS_COMPRESSED_READ  (26),
		.IN_PKT_BURSTWRAP_H            (37),
		.IN_PKT_BURSTWRAP_L            (35),
		.IN_PKT_BURST_SIZE_H           (40),
		.IN_PKT_BURST_SIZE_L           (38),
		.IN_PKT_RESPONSE_STATUS_H      (64),
		.IN_PKT_RESPONSE_STATUS_L      (63),
		.IN_PKT_TRANS_EXCLUSIVE        (31),
		.IN_PKT_BURST_TYPE_H           (42),
		.IN_PKT_BURST_TYPE_L           (41),
		.IN_ST_DATA_W                  (65),
		.OUT_PKT_ADDR_H                (52),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (61),
		.OUT_PKT_BYTE_CNT_L            (59),
		.OUT_PKT_TRANS_COMPRESSED_READ (53),
		.OUT_PKT_BURST_SIZE_H          (67),
		.OUT_PKT_BURST_SIZE_L          (65),
		.OUT_PKT_RESPONSE_STATUS_H     (91),
		.OUT_PKT_RESPONSE_STATUS_L     (90),
		.OUT_PKT_TRANS_EXCLUSIVE       (58),
		.OUT_PKT_BURST_TYPE_H          (69),
		.OUT_PKT_BURST_TYPE_L          (68),
		.OUT_ST_DATA_W                 (92),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_004_src_valid),             //      sink.valid
		.in_channel           (id_router_004_src_channel),           //          .channel
		.in_startofpacket     (id_router_004_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_004_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_004_src_ready),             //          .ready
		.in_data              (id_router_004_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (52),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (61),
		.IN_PKT_BYTE_CNT_L             (59),
		.IN_PKT_TRANS_COMPRESSED_READ  (53),
		.IN_PKT_BURSTWRAP_H            (64),
		.IN_PKT_BURSTWRAP_L            (62),
		.IN_PKT_BURST_SIZE_H           (67),
		.IN_PKT_BURST_SIZE_L           (65),
		.IN_PKT_RESPONSE_STATUS_H      (91),
		.IN_PKT_RESPONSE_STATUS_L      (90),
		.IN_PKT_TRANS_EXCLUSIVE        (58),
		.IN_PKT_BURST_TYPE_H           (69),
		.IN_PKT_BURST_TYPE_L           (68),
		.IN_ST_DATA_W                  (92),
		.OUT_PKT_ADDR_H                (25),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (34),
		.OUT_PKT_BYTE_CNT_L            (32),
		.OUT_PKT_TRANS_COMPRESSED_READ (26),
		.OUT_PKT_BURST_SIZE_H          (40),
		.OUT_PKT_BURST_SIZE_L          (38),
		.OUT_PKT_RESPONSE_STATUS_H     (64),
		.OUT_PKT_RESPONSE_STATUS_L     (63),
		.OUT_PKT_TRANS_EXCLUSIVE       (31),
		.OUT_PKT_BURST_TYPE_H          (42),
		.OUT_PKT_BURST_TYPE_L          (41),
		.OUT_ST_DATA_W                 (65),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_mux_006_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_006_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_006_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_006_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_006_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_006_src_data),           //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (25),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (34),
		.IN_PKT_BYTE_CNT_L             (32),
		.IN_PKT_TRANS_COMPRESSED_READ  (26),
		.IN_PKT_BURSTWRAP_H            (37),
		.IN_PKT_BURSTWRAP_L            (35),
		.IN_PKT_BURST_SIZE_H           (40),
		.IN_PKT_BURST_SIZE_L           (38),
		.IN_PKT_RESPONSE_STATUS_H      (64),
		.IN_PKT_RESPONSE_STATUS_L      (63),
		.IN_PKT_TRANS_EXCLUSIVE        (31),
		.IN_PKT_BURST_TYPE_H           (42),
		.IN_PKT_BURST_TYPE_L           (41),
		.IN_ST_DATA_W                  (65),
		.OUT_PKT_ADDR_H                (52),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (61),
		.OUT_PKT_BYTE_CNT_L            (59),
		.OUT_PKT_TRANS_COMPRESSED_READ (53),
		.OUT_PKT_BURST_SIZE_H          (67),
		.OUT_PKT_BURST_SIZE_L          (65),
		.OUT_PKT_RESPONSE_STATUS_H     (91),
		.OUT_PKT_RESPONSE_STATUS_L     (90),
		.OUT_PKT_TRANS_EXCLUSIVE       (58),
		.OUT_PKT_BURST_TYPE_H          (69),
		.OUT_PKT_BURST_TYPE_L          (68),
		.OUT_ST_DATA_W                 (92),
		.ST_CHANNEL_W                  (9),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_003 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_006_src_valid),             //      sink.valid
		.in_channel           (id_router_006_src_channel),           //          .channel
		.in_startofpacket     (id_router_006_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_006_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_006_src_ready),             //          .ready
		.in_data              (id_router_006_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

endmodule
